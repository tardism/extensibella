grammar extensibella:fromAbella;

exports extensibella:fromAbella:abstractSyntax;
exports extensibella:fromAbella:concreteSyntax;
