grammar extensibella:common;

exports extensibella:common:abstractSyntax;
exports extensibella:common:concreteSyntax;
