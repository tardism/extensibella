grammar extensibella:toAbella:abstractSyntax;

imports extensibella:common:abstractSyntax;
