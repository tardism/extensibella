grammar extensibella:outerfaceFile;

exports extensibella:outerfaceFile:concreteSyntax;
exports extensibella:outerfaceFile:abstractSyntax;
