grammar extensibella:fromAbella:abstractSyntax;

