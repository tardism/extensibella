grammar extensibella:toAbella;

exports extensibella:toAbella:abstractSyntax;
exports extensibella:toAbella:concreteSyntax;
