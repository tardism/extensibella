grammar extensibella:interfaceFile;

exports extensibella:interfaceFile:concreteSyntax;
exports extensibella:interfaceFile:abstractSyntax;
